-------------------------------------------------------------------------
-- Joseph Zambreno
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- invg.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of a 1-input NOT 
-- gate.
--
--
-- NOTES:
-- 8/19/16 by JAZ::Design created.
-- 1/16/19 by H3::Changed name to avoid name conflict with Quartus 
--         primitives.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
entity decoder_5to32 is
  port(i_A          : in std_logic_vector(4 downto 0);
       Enable	    : in std_logic;
       o_F          : out std_logic_vector(31 downto 0));
end decoder_5to32;

architecture dataflow of decoder_5to32 is
signal concat : std_logic_vector(5 downto 0);
begin
concat <= i_A & Enable;
	 with concat select o_F <=
		"00000000000000000000000000000001" when "000001",
		"00000000000000000000000000000010" when "000011",
		"00000000000000000000000000000100" when "000101",
		"00000000000000000000000000001000" when "000111",
		"00000000000000000000000000010000" when "001001",
		"00000000000000000000000000100000" when "001011",
		"00000000000000000000000001000000" when "001101",
		"00000000000000000000000010000000" when "001111",
		"00000000000000000000000100000000" when "010001",
		"00000000000000000000001000000000" when "010011",
		"00000000000000000000010000000000" when "010101",
		"00000000000000000000100000000000" when "010111",
		"00000000000000000001000000000000" when "011001",
		"00000000000000000010000000000000" when "011011",
		"00000000000000000100000000000000" when "011101",
		"00000000000000001000000000000000" when "011111",
		"00000000000000010000000000000000" when "100001",
		"00000000000000100000000000000000" when "100011",
		"00000000000001000000000000000000" when "100101",
		"00000000000010000000000000000000" when "100111",
		"00000000000100000000000000000000" when "101001",
		"00000000001000000000000000000000" when "101011",
		"00000000010000000000000000000000" when "101101",
		"00000000100000000000000000000000" when "101111",
		"00000001000000000000000000000000" when "110001",
		"00000010000000000000000000000000" when "110011",
		"00000100000000000000000000000000" when "110101",
		"00001000000000000000000000000000" when "110111",
		"00010000000000000000000000000000" when "111001",
		"00100000000000000000000000000000" when "111011",
		"01000000000000000000000000000000" when "111101",
		"10000000000000000000000000000000" when "111111",
		"00000000000000000000000000000000" when others;
end dataflow;