-------------------------------------------------------------------------
-- Henry Duwe
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- MIPS_Processor.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains a skeleton of a MIPS_Processor  
-- implementation.

-- 01/29/2019 by H3::Design created.
-------------------------------------------------------------------------


library IEEE;
use IEEE.std_logic_1164.all;


entity MIPS_Processor is
  generic(N : integer := 32);
  port(iCLK            : in std_logic;
       iRST            : in std_logic;
       iInstLd         : in std_logic;
       iInstAddr       : in std_logic_vector(N-1 downto 0);
       iInstExt        : in std_logic_vector(N-1 downto 0);
       oALUOut         : out std_logic_vector(N-1 downto 0)); -- TODO: Hook this up to the output of the ALU. It is important for synthesis that you have this output that can effectively be impacted by all other components so they are not optimized away.

end  MIPS_Processor;


architecture structure of MIPS_Processor is

  -- Required data memory signals
  signal s_DMemWr       : std_logic; -- TODO: use this signal as the final active high data memory write enable signal
  signal s_DMemAddr     : std_logic_vector(N-1 downto 0); -- TODO: use this signal as the final data memory address input
  signal s_DMemData     : std_logic_vector(N-1 downto 0); -- TODO: use this signal as the final data memory data input
  signal s_DMemOut      : std_logic_vector(N-1 downto 0); -- TODO: use this signal as the data memory output
 
  -- Required register file signals 
  signal s_RegWr        : std_logic; -- TODO: use this signal as the final active high write enable input to the register file
  signal s_RegWrAddr    : std_logic_vector(4 downto 0); -- TODO: use this signal as the final destination register address input
  signal s_RegWrData    : std_logic_vector(N-1 downto 0); -- TODO: use this signal as the final data memory data input

  -- Required instruction memory signals
  signal s_IMemAddr     : std_logic_vector(N-1 downto 0); -- Do not assign this signal, assign to s_NextInstAddr instead
  signal s_NextInstAddr : std_logic_vector(N-1 downto 0); -- TODO: use this signal as your intended final instruction memory address input.
  signal s_Inst         : std_logic_vector(N-1 downto 0); -- TODO: use this signal as the instruction signal 

  -- Required halt signal -- for simulation
  signal v0             : std_logic_vector(N-1 downto 0); -- TODO: should be assigned to the output of register 2, used to implement the halt SYSCALL
  signal s_Halt         : std_logic;  -- TODO: this signal indicates to the simulation that intended program execution has completed. This case happens when the syscall instruction is observed and the V0 register is at 0x0000000A. This signal is active high and should only be asserted after the last register and memory writes before the syscall are guaranteed to be completed.

  component mem is
    generic(ADDR_WIDTH : integer;
            DATA_WIDTH : integer);
    port(
          clk          : in std_logic;
          addr         : in std_logic_vector((ADDR_WIDTH-1) downto 0);
          data         : in std_logic_vector((DATA_WIDTH-1) downto 0);
          we           : in std_logic := '1';
          q            : out std_logic_vector((DATA_WIDTH -1) downto 0));
    end component;

  -- TODO: You may add any additional signals or components your implementation 
  --       requires below this comment
  
  component register_file
port(i_CLK          : in std_logic;     -- Clock input
     i_Res	    : in std_logic;   -- Reset
     i_We           : in std_logic_vector(4 downto 0);	-- Write address input
     i_Re1          : in std_logic_vector(4 downto 0);  --Read enable input
     i_Re2          : in std_logic_vector(4 downto 0);	--Read enable input
     i_D            : in std_logic_vector(31 downto 0);	-- Data value input
     i_WrEn	    : in std_logic;
     out1           : out std_logic_vector(31 downto 0);   -- Data value output   
     out2           : out std_logic_vector(31 downto 0);
     v0             : out std_logic_vector(31 downto 0));   -- Data value output
  end component;
component ALUSHIFT
  port(i_A : in std_logic_vector(31 downto 0);
	i_B : in std_logic_vector(31 downto 0);
	i_Im : in std_logic_vector(31 downto 0);
	i_Binv : in std_logic;
	ALUsrc : in std_logic;
	i_Op : in std_logic_vector(5 downto 0);
	i_Shift : in std_logic_vector(4 downto 0);
	o_Out : out std_logic_vector(31 downto 0);
        o_Zero : out std_logic);				    
end component;


component mux
port(i_s	    : in std_logic;
       i_A          : in std_logic_vector(31 downto 0);
       i_B	    : in std_logic_vector(31 downto 0);
       o_y         : out std_logic_vector(31 downto 0));
end component;

component signExtend
port(i_A : in std_logic_vector(15 downto 0);
     i_Sel : in std_logic;
     o_Out : out std_logic_vector(31 downto  0));
end component;

component PC is
  port(i_CLK        : in std_logic;     -- Clock input
       i_RST        : in std_logic;     -- Reset input
       i_WE         : in std_logic;     -- Write enable input
       i_D          : in std_logic_vector(31 downto 0);     -- Data value input
       o_Q          : out std_logic_vector(31 downto 0));   -- Data value output
end component;

component full_adder is
port(i_A          : in std_logic_vector(31 downto 0);
       i_B          : in std_logic_vector(31 downto 0);
       o_S          : out std_logic_vector(31 downto 0);
       i_C          : in std_logic;
       o_C          : out std_logic);

end component;

component mux5bit is
generic(N : integer := 5);
  port(sel	    : in std_logic;
       i_A          : in std_logic_vector(N-1 downto 0);
       i_B	    : in std_logic_vector(N-1 downto 0);
       o_F          : out std_logic_vector(N-1 downto 0));

end component;

component IFID is
  port(i_CLK        : in std_logic;     -- Clock input
       iWrEn        : in std_logic;	-- Write enable input
       iRst         : in std_logic;     -- Reset input
       iInstruction : in std_logic_vector(31 downto 0);     -- Data value input
       iPC4         : in std_logic_vector(31 downto 0);
       o_Q          : out std_logic_vector(63 downto 0));   -- Data value output
end component;
component controlModule is
  port(opCode       : in std_logic_vector(5 downto 0);
       functCode    : in std_logic_vector(5 downto 0);
       RegDst       : out std_logic;
       MemToReg	    : out std_logic;
       ALUOp	    : out std_logic_vector(5 downto 0);
       MemWrite     : out std_logic;
       ALUSrc       : out std_logic;
       RegWrite     : out std_logic;
       BInvert      : out std_logic;
       SelExt	    : out std_logic;
       SelLui	    : out std_logic;
       SelShift     : out std_logic;
       SelBranch    : out std_logic;
       branch       : out std_logic;
       jump         : out std_logic;
       jal	    : out std_logic;
       jr           : out std_logic);

end component;

component shift2 is
  port(i_A   : in std_logic_vector(31 downto 0);
       o_Y : out std_logic_vector(31 downto 0));
end component;

component mux1bit is
  port(sel	    : in std_logic;
       i_A          : in std_logic;
       i_B	    : in std_logic;
       o_F          : out std_logic);
end component;

component andg2 is
  port(i_A          : in std_logic;
       i_B          : in std_logic;
       o_F          : out std_logic);
end component;

component invg is
  port(i_A          : in std_logic;
       o_F          : out std_logic);
end component;

component padder is
  port(i_A   : in std_logic_vector(15 downto 0);
       o_Y : out std_logic_vector(31 downto 0));
end component;

component jumpShift2 is
  port(i_A   : in std_logic_vector(25 downto 0);
       o_Y   : out std_logic_vector(27 downto 0));

end component;
component Compare is
  port(i_A : in std_logic_vector(31 downto 0);
       i_B : in std_logic_vector(31 downto 0);
       o_Q : out std_logic);

end component;

component IDEX is
  port(i_CLK        : in std_logic;-- Clock input
       iRst         : in std_logic;
       iWrEn        : in std_logic;	-- Write enable input
       iRegDst      : in std_logic;
       iMemToReg    : in std_logic;
       iALUOp	    : in std_logic_vector(5 downto 0);
       iMemWrite    : in std_logic;
       iALUSrc      : in std_logic;
       iRegWrite    : in std_logic;
       iBInvert     : in std_logic;
       iSelExt	    : in std_logic;
       iSelLui	    : in std_logic;
       iSelShift    : in std_logic;
       iPC4         : in std_logic_vector(31 downto 0);
       i_A	    : in std_logic_vector(31 downto 0);
       i_B 	    : in std_logic_vector(31 downto 0);
       i_Im	    : in std_logic_vector(31 downto 0);
       i_Rt         : in std_logic_vector(4 downto 0);
       i_Rd         : in std_logic_vector(4 downto 0);
       oRegDst      : out std_logic;
       oMemToReg    : out std_logic;
       oALUOp	    : out std_logic_vector(5 downto 0);
       oMemWrite    : out std_logic;
       oALUSrc      : out std_logic;
       oRegWrite    : out std_logic;
       oBinvert     : out std_logic;
       oSelExt	    : out std_logic;
       oSelLui	    : out std_logic;
       oSelShift    : out std_logic;
       oPC4         : out std_logic_vector(31 downto 0);
       o_A	    : out std_logic_vector(31 downto 0);
       o_B          : out std_logic_vector(31 downto 0);
       o_Im	    : out std_logic_vector(31 downto 0);
       o_Rt         : out std_logic_vector(4 downto 0);
       o_Rd         : out std_logic_vector(4 downto 0));
      

end component;
component EXMEM is
  port(i_CLK        : in std_logic;-- Clock input
       iRst         : in std_logic;
       iWrEn        : in std_logic;	-- Write enable input
       iMemToReg    : in std_logic;
       iMemWrite    : in std_logic;
       iRegWrite    : in std_logic;
       iSelLui	    : in std_logic;
       i_B 	    : in std_logic_vector(31 downto 0);
       i_RealRd     : in std_logic_vector(4 downto 0);
       i_ALUOut     : in std_logic_vector(31 downto 0);
       i_Inst       : in std_logic_vector(15 downto 0);
       oMemToReg    : out std_logic;
       oMemWrite    : out std_logic;
       oRegWrite    : out std_logic;
       oSelLui	    : out std_logic;
       o_B 	    : out std_logic_vector(31 downto 0);
       o_RealRd     : out std_logic_vector(4 downto 0);
       o_ALUOut     : out std_logic_vector(31 downto 0);
       o_Inst       : out std_logic_vector(15 downto 0));
      

end component;

component MEMWB is
  port(i_CLK        : in std_logic;-- Clock input
       iRst         : in std_logic;
       iWrEn        : in std_logic;	-- Write enable input
       iMemToReg    : in std_logic;
       iRegWrite    : in std_logic;
       iSelLui	    : in std_logic;
       iDMemOut     : in std_logic_vector(31 downto 0);
       iDMemAddr    : in std_logic_vector(31 downto 0);
       iRealRd      : in std_logic_vector(4 downto 0);
       iIm          : in std_logic_vector(15 downto 0);
       oMemToReg    : out std_logic;
       oRegWrite    : out std_logic;
       oSelLui	    : out std_logic;
       oDMemOut     : out std_logic_vector(31 downto 0);
       oDMemAddr    : out std_logic_vector(31 downto 0);
       oIm          : out std_logic_vector(15 downto 0);
       oRealRd      : out std_logic_vector(4 downto 0));
end component;

signal s_A1, s_Im,wb_DMemOut, wb_DMemAddr,s_PCNEW, s_MemLui, s_branchShift2, s_branchAddr, s_PCFinal, s_padLUI, s_PCBranch, s_JumpAdr, s_RegData, s_PCBranchJump, id_DMemData, ex_Im, ex_A, ex_B, mem_ALUOut, ex_DMemAddr : std_logic_vector(31 downto 0);
signal s_Zero,wb_MemToReg,wb_RegWrite, s_RegDst, s_MemToReg,wb_SelLui, s_ALUSrc, s_BInvert, s_SelExt, s_SelLui, s_ShiftVar, s_SelBranch, s_branch, s_isBranch, s_beqAND, s_bneAND, s_notZero, s_jump, s_jal, s_Jr , id_RegWr, id_DMemWr, ex_RegDst, ex_MemToReg, ex_MemWrite, ex_ALUSrc, ex_RegWrite, ex_BInvert, ex_SelExt, ex_SelLui, ex_SelShift, mem_MemToReg, mem_MemWrite, mem_RegWrite, mem_SelLui, mem_B : std_logic;
signal s_ALUOp, ex_ALUOp : std_logic_vector(5 downto 0);
signal mem_Inst,wb_Im : std_logic_vector(15 downto 0);
signal s_ShiftAm,wb_RealRD,mem_RealRD, s_RSRT, ex_Rt, ex_Rd : std_logic_vector(4 downto 0);
signal s_jumpShift2: std_logic_vector(27 downto 0);
signal  s_IFIDOut : std_logic_vector(63 downto 0);







begin

  -- TODO: This is required to be your final input to your instruction memory. This provides a feasible method to externally load the memory module which means that the synthesis tool must assume it knows nothing about the values stored in the instruction memory. If this is not included, much, if not all of the design is optimized out because the synthesis tool will believe the memory to be all zeros.
  with iInstLd select
    s_IMemAddr <= s_NextInstAddr when '0',
      iInstAddr when others;


  IMem: mem
    generic map(ADDR_WIDTH => 10,
                DATA_WIDTH => N)
    port map(clk  => iCLK,
             addr => s_IMemAddr(11 downto 2),
             data => iInstExt,
             we   => iInstLd,
             q    => s_Inst);
  
  DMem: mem
    generic map(ADDR_WIDTH => 10,
                DATA_WIDTH => N)
    port map(clk  => iCLK,
             addr => s_DMemAddr(11 downto 2),
             data => s_DMemData,
             we   => s_DMemWr,
             q    => s_DMemOut);

  s_Halt <='1' when (s_Inst(31 downto 26) = "000000") and (s_Inst(5 downto 0) = "001100") and (v0 = "00000000000000000000000000001010") else '0';

  -- TODO: Implement the rest of your processor below this comment! 
  g_PC: PC
	port map(i_CLK => iCLK,
		 i_RST => iRST,
		 i_WE => '1',
		 i_D => s_PCFinal,
		 o_Q => s_NextInstAddr);
 adder: full_adder
	port map(i_A => s_NextInstAddr,
		 i_B => x"00000004",
		 o_S => s_PCNEW,
		 i_C => '0',
		 o_C => open);
 a_IFID: IFID
	port map(i_CLK => iCLK,
       		iWrEn => '1',
      		iRst => '0',
      		iInstruction => s_Inst,
       		iPC4 => s_PCNEW,
       		o_Q => s_IFIDOut);

control: controlModule
	port map(opCode => s_IFIDOut(31 downto 26),
		 functCode => s_IFIDOut(5 downto 0),
		 RegDst => s_RegDst,
		 MemToReg => s_MemToReg,
		 ALUOp => s_ALUOp,
		 MemWrite => id_DMemWr,
		 ALUSrc => s_ALUSrc,
		 RegWrite => id_RegWr,
		 BInvert => s_BInvert,
		 SelExt => s_SelExt,
		 SelLui => s_SelLui,
		 SelShift => s_ShiftVar,
		 SelBranch => s_SelBranch,
		 branch  => s_branch,
                 jump => s_jump,
		 jal => s_jal,
		 jr  => s_Jr);


extender: signExtend
	port map(i_A => s_IFIDOut(15 downto 0),
    		 i_Sel => s_SelExt,
    		 o_Out => s_Im);

bZero: compare
	port map(i_A => s_A1,
		 i_B => id_DMemData,
	         o_Q => s_Zero);

muxPC: mux
	port map(i_s => s_jal,
		 i_A => s_RegData,
		 i_B => s_PCNew,
	         o_y => s_RegWrData);

branchShift2: shift2
  	port map(i_A => s_Im,
                 o_Y => s_branchShift2);

muxSelBranch: mux1bit
	port map(sel => s_SelBranch,
	         i_A => s_bneAND,
	         i_B => s_beqAND,
	         o_F => s_isBranch);

BranchAdder: full_adder
	port map(i_A => s_PCNEW,
		 i_B => s_branchShift2,
		 o_S => s_branchAddr,
		 i_C => '0',
		 o_C => open);		 

muxAddr: mux
	port map(i_s => s_isBranch,
		 i_A => s_PCNEW,
	         i_B => s_branchAddr,
	         o_y => s_PCBranch);

beqAnd: andg2
	port map(i_A => s_branch,
                 i_B => s_Zero,
		 o_F => s_beqAND);

nZero: invg
	port map(i_A => s_Zero,
                 o_F => s_notZero);

bneAND: andg2
	port map(i_A => s_branch,
                 i_B => s_notZero,
                 o_F => s_bneAND);

g_jumpShift2: jumpShift2
  	port map(i_A => s_IFIDOut(25 downto 0),
                 o_Y => s_jumpShift2);

s_JumpAdr <= s_PCNEW(31 downto 28) & s_jumpShift2;

muxJump: mux
	port map(i_s => s_jump,
		 i_A => s_PCBranch,
	         i_B => s_JumpAdr,
	         o_y => s_PCBranchJump);
muxWrAddr: mux5bit
	port map(sel => s_jal,
		 i_A => wb_RealRD,
		 i_B => "11111",
		 o_F => s_RegWrAddr);
muxJR: mux
	port map(i_s => s_Jr,
		 i_A => s_PCBranchJump,
		 i_B => s_A1,
		 o_Y => s_PCFINAL);

reg: register_file
	port map(i_CLK => iCLK,
     		i_Res => iRST,	    
     		i_We  => s_RegWrAddr,   
     		i_Re1  => s_IFIDOut(25 downto 21),    
     		i_Re2   => s_IFIDOut(20 downto 16),   
     		i_D      => s_RegWrData,  
     		i_WrEn	 =>  s_RegWrite,
     		out1     => s_A1,
	        out2 => id_DMemData,
	        v0 => v0);

aIDEX: IDEX
 port map(i_CLK=> iCLK,
       iRst => '0',
       iWrEn => '1',
       iRegDst => s_RegDst,
       iMemToReg => s_MemtoReg,
       iALUOp => s_ALUOp,
       iMemWrite => id_DMemWr,
       iALUSrc => s_ALUSrc,
       iRegWrite => id_RegWr,
       iBInvert =>s_BInvert,
       iSelExt => s_SelExt,
       iSelLui => s_SelLui,
       iSelShift => s_ShiftVar,
       iPC4 => s_PCNEW,
       i_A => s_A1,
       i_B => id_DMemData,
       i_Im => s_Im,
       i_Rt => s_IFIDOut(20 downto 16),
       i_Rd  => s_IFIDOut(15 downto 11),
       oRegDst => ex_RegDst,
       oMemToReg => ex_MemToReg,
       oALUOp => ex_ALUOp,
       oMemWrite => ex_MemWrite,
       oALUSrc => ex_ALUSrc,
       oRegWrite => ex_RegWrite,
       oBinvert => ex_BInvert,
       oSelExt => ex_SelExt,
       oSelLui	=> ex_SelLui,
       oSelShift => ex_SelShift,
       oPC4 => open,
       o_A => ex_A,
       o_B => ex_B,
       o_Im => ex_Im,
       o_Rt => ex_Rt,
       o_Rd => ex_Rd);

mux1: mux5bit
	port map(sel => ex_RegDst,
		 i_A => ex_Rt,
		 i_B => ex_Rd,
		 o_F => s_RSRT);
mux2: mux5bit
	port map(sel =>	ex_SelShift,
		 i_A => ex_Rt,
		 i_B => s_A1(4 downto 0),
		 o_F => s_ShiftAm);
alu: ALUSHIFT
	port map(i_A => ex_A,
		i_B => ex_B,
		i_Im => ex_Im,
		i_Binv => ex_BInvert,
		ALUsrc => ex_ALUSrc,
		i_Op => ex_ALUOp,
		i_Shift => s_ShiftAm,
		o_Out => ex_DMemAddr,
        	o_Zero => open);

aEXMEM: EXMEM
port map(i_CLK => iCLK,
       iRst => '0',
       iWrEn => '1',
       iMemToReg => ex_MemToReg,
       iMemWrite => ex_MemWrite,
       iRegWrite => ex_RegWrite, --Ask ta about reg write for jal
       iSelLui => ex_SelLui,
       i_B => ex_B,
       i_RealRd => s_RSRT,
       i_ALUOut => ex_DmemAddr,
       i_Inst  => ex_Im(15 downto 0),
       oMemToReg => mem_MemToReg,
       oMemWrite => s_DmemWr,
       oRegWrite => mem_RegWrite,
       oSelLui	 => mem_SelLui,
       o_B 	 => s_DmemData,
       o_RealRd  => mem_RealRD,
       o_ALUOut  => s_DmemAddr,
       o_Inst    => mem_Inst);


aMEMWB : MEMWB
 port map(i_CLK => iCLK,
       iRst => '0',
       iWrEn => '1',
       iMemToReg => mem_MemToReg,
       iRegWrite => mem_RegWrite,
       iSelLui	 => mem_SelLui,
       iDMemOut  => s_DMemOut,
       iDMemAddr  => s_DmemAddr,
       iRealRd    => mem_RealRD,
       iIm        => mem_Inst,
       oMemToReg  => wb_MemToReg,
       oRegWrite  => s_RegWrite,
       oSelLui	  => wb_SelLui,
       oDMemOut   => wb_DMemOut,
       oDMemAddr  => wb_DMemAddr,
       oIm        => wb_Im,
       oRealRd    => wb_RealRD);

muxAluMem: mux
	port map(i_s => wb_MemToReg,
      		 i_A => wb_DMemAddr,
       		 i_B => wb_DmemOut,
       		 o_y => s_MemLui);
padLUI: padder
	port map(i_A => wb_Im,
		 o_Y => s_padLUI);

muxLUI: mux
	port map(i_s => wb_SelLui,
		 i_A => s_MemLui,
		 i_B => s_padLUI,
	         o_y => s_RegData);
end structure;
