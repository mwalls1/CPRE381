-------------------------------------------------------------------------
-- Joseph Zambreno
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- dff.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of an edge-triggered
-- flip-flop with parallel access and reset.
--
--
-- NOTES:
-- 8/19/16 by JAZ::Design created.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity add_sub_reg is
  port(i_CLK        : in std_logic;     -- Clock input
       i_Res        : in std_logic;	-- Reset input
       i_WrEn       : in std_logic;     -- Global write enable
       i_We         : in std_logic_vector(4 downto 0);-- Write address input
       i_Re1        : in std_logic_vector(4 downto 0);--Read Address input
       i_Re2        : in std_logic_vector(4 downto 0);--Read Address input
       i_Im         : in std_logic_vector(31 downto 0);--Immediate input
       i_Add_Sub    : in std_logic;
       i_ALUSRc	    : in std_logic);					    

end add_sub_reg;

architecture structure of add_sub_reg is
component register_file
port(i_CLK          : in std_logic;     -- Clock input
     i_Res	    : in std_logic;   -- Reset
     i_We           : in std_logic_vector(4 downto 0);	-- Write enable input
     i_Re1          : in std_logic_vector(4 downto 0);  --Read enable input
     i_Re2          : in std_logic_vector(4 downto 0);	--Read enable input
     i_D            : in std_logic_vector(31 downto 0);	-- Data value input
     i_WrEn	    : in std_logic;
     out1           : out std_logic_vector(31 downto 0);   -- Data value output   
     out2           : out std_logic_vector(31 downto 0));   -- Data value output
  end component;
component add_sub
port(nAdd_Sub			    : in std_logic;
       ALUSrc			    : in std_logic;
       iA 		            : in std_logic_vector(31 downto 0);
       iB 		            : in std_logic_vector(31 downto 0);
       iIm			    : in std_logic_vector(31 downto 0);
       sum 		            : out std_logic_vector(31 downto 0);
       Co			    : out std_logic);
end component;

signal s_Sum, s_A1, s_A2 : std_logic_vector(31 downto 0);

begin

g_r1 : register_file
	port MAP(i_CLK => i_CLK,
		i_Res => i_Res,
		i_We => i_We,
		i_Re1 => i_Re1,
		i_Re2 => i_Re2,
		i_D => s_Sum,
		i_WrEn => i_WrEn,
		out1 => s_A1,
		out2 => s_A2);
g_add1 : add_sub
	port MAP(nAdd_Sub => i_Add_Sub,
		ALUSrc => i_ALUSRc,
		iA => s_A1,
		iB => s_A2,
		iIm => i_Im,
		sum => s_Sum,
		Co => OPEN);
end structure;