library IEEE;
use IEEE.std_logic_1164.all;

entity Concatenate is
port(i_X  : in std_logic_vector(31 downto 0);
     i_Am : in integer;
     o_Y  : out std_logic_vector(31 downto 0));
end Concatenate;

architecture dataflow of Concatenate is

signal temp : std_logic_vector (31 downto 0);

begin
  temp <= i_X (30 downto 0) & '0';

   G: for i in 0 to i_Am generate
	temp <= temp(30 downto 0) & '0';
   end generate;

o_Y <= temp;
end dataflow;